`timescale 1ns / 1ps

module GCD(
    input [7:0] X,Y,
	 input clk,
    output [7:0] GCD
    );

always @(negedge clk)
begin
	
end

endmodule
